// SPDX-License-Identifier: AGPL-3.0-Only
/*
 * Copyright (C) 2022 Sean Anderson <seanga2@gmail.com>
 */

`ifndef COMMON_VH
`define COMMON_VH

`default_nettype none
`timescale 1ns/1ns

`endif /* COMMON_VH */
