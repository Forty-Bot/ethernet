`ifndef IO_VH
`define IO_VH

`define PIN_INPUT_REGISTERED		6'b000000
`define PIN_INPUT_UNREGISTERED		6'b000001
`define PIN_INPUT_LATCH			6'b000010
`define PIN_INPUT_DDR			6'b000000

`define PIN_OUTPUT_NEVER		6'b000000
`define PIN_OUTPUT_ALWAYS		6'b010000
`define PIN_OUTPUT_ENABLE		6'b100000
`define PIN_OUTPUT_ENABLE_REGISTERED	6'b110000

`define PIN_OUTPUT_DDR			6'b000000
`define PIN_OUTPUT_REGISTERED		6'b000100
`define PIN_OUTPUT_UNREGISTERED		6'b001000
`define PIN_OUTPUT_REGISTERED_INVERTED	6'b001100

`endif /* IO_VH */
